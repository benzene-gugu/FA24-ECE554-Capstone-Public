00
c0
00
c7
00
f5
07
f5
17
d7
5f
00
07
07
f6
06
00
a7
00
00
07
87
07
00
47
f5
00
01
81
21
11
91
05
40
04
f9
84
94
5f
95
a4
09
c1
81
41
01
01
00
01
fa
11
81
91
21
31
41
51
61
f7
00
e7
00
07
c4
f4
04
00
00
00
f4
07
1f
04
07
37
f7
50
19
00
c0
35
00
f4
10
f4
00
07
00
e7
df
44
f9
09
10
5f
00
00
00
00
c9
04
89
09
09
0a
04
94
40
9a
99
04
00
fa
f7
00
d7
e7
00
07
00
07
00
04
10
a0
30
44
1f
35
55
00
f4
df
41
5f
c1
df
00
00
41
f4
81
5f
81
25
a0
5f
04
9f
c1
5f
a9
9b
ab
14
1f
04
9f
41
1f
41
07
1f
00
07
15
15
85
f7
a7
f7
00
00
47
a5
15
00
00
47
35
35
00
00
47
65
35
00
00
07
15
95
f7
a7
f7
00
01
81
91
21
11
05
05
06
5f
05
5f
05
00
00
e7
00
00
87
87
1f
85
00
00
e7
10
df
df
05
1f
5f
85
00
00
e7
00
00
c7
87
1f
05
00
00
e7
c1
81
41
01
01
00
f9
06
17
d7
5f
07
f4
17
c6
df
01
f0
10
11
f1
1f
c1
81
40
1f
00
9f
d1
e1
f1
c1
07
87
e7
a7
01
00
01
21
11
81
91
31
46
00
27
c1
81
00
00
e7
41
01
c1
01
00
00
30
e7
05
e7
85
05
05
85
b7
05
10
06
e7
00
5f
5f
05
5f
05
00
00
e7
00
00
87
27
1f
25
00
00
e7
10
df
df
05
1f
5f
25
00
00
e7
00
c7
c7
e4
07
e4
07
e4
07
e4
00
97
1f
05
00
07
00
e7
81
c1
41
01
c1
00
01
5f
f9
06
17
d7
9f
07
e4
17
c6
1f
