37
ef
93
63
67
33
83
33
93
23
6f
37
83
93
93
e3
b7
23
67
37
83
93
e3
b7
03
13
67
13
23
23
23
23
13
13
83
13
93
23
ef
33
23
e3
83
03
83
03
13
67
13
b7
23
23
23
23
23
23
23
23
93
73
e3
b7
03
13
13
63
b7
93
37
23
83
b7
93
93
93
23
13
93
13
ef
63
93
23
93
63
b7
93
13
23
6f
23
13
e3
13
6f
37
93
13
37
13
93
63
93
93
13
13
33
ef
33
b3
e3
f3
b7
93
73
33
e3
b7
23
93
e7
37
13
13
93
93
23
ef
63
e3
93
23
ef
13
ef
13
ef
93
13
83
63
13
ef
03
33
33
ef
23
6f
03
ef
33
33
23
93
6f
23
ef
13
ef
83
e7
6f
37
83
13
13
13
93
b3
23
67
b7
03
13
13
67
b7
03
13
13
67
b7
03
13
13
67
37
83
13
13
93
b3
23
67
13
23
23
23
23
13
93
13
ef
e3
ef
63
b7
13
23
37
93
13
63
ef
63
b7
13
23
13
ef
ef
e3
ef
ef
63
b7
13
23
37
93
13
63
ef
63
b7
13
23
83
03
83
03
13
67
b3
83
93
23
6f
03
b3
93
23
6f
13
93
13
23
23
ef
93
13
13
ef
13
ef
83
03
03
83
93
13
b3
33
13
67
13
23
23
23
23
23
13
b7
63
83
03
b7
13
23
83
03
83
13
67
93
13
23
13
a3
13
93
93
93
33
13
13
93
23
93
ef
ef
e3
ef
63
b7
13
23
37
93
13
63
ef
63
b7
13
23
13
ef
ef
e3
ef
ef
63
b7
13
23
b7
03
93
23
03
23
03
23
03
23
13
63
ef
63
b7
93
13
23
03
83
83
03
83
13
13
6f
b3
83
93
23
6f
03
b3
13
23
6f
