04
0b
00
00
00
00
00
00
00
00
fe
10
00
01
0f
fe
10
00
00
10
00
01
fe
10
00
0f
00
ff
00
01
00
00
00
00
00
ff
00
00
fb
00
00
fe
00
00
00
00
01
00
fd
02
02
02
02
03
01
01
01
01
07
c0
fe
10
02
00
0f
0e
10
20
11
00
00
00
01
f0
00
00
00
90
10
2b
03
20
00
00
02
10
01
10
00
ff
01
ff
fc
00
fd
00
00
00
01
ff
00
00
00
00
00
00
40
2a
00
00
fc
c0
02
07
c0
40
fe
10
00
00
00
10
01
00
06
07
01
e5
07
ff
20
00
e1
00
e5
00
e4
00
00
00
02
00
e3
00
41
00
de
00
fa
00
df
00
00
00
00
fc
00
db
00
df
00
00
f7
11
00
00
00
00
ef
00
00
00
11
00
01
00
00
11
00
01
01
00
11
00
00
01
00
11
00
00
00
df
00
00
00
ff
00
00
01
00
00
00
00
f8
fe
fa
00
10
10
00
11
00
00
06
f8
00
10
10
00
00
f7
f3
fe
f7
f4
00
10
10
00
11
00
00
04
f2
00
10
10
00
00
00
00
00
01
00
00
00
00
00
f7
00
00
00
00
fa
fe
09
00
00
00
e8
00
00
00
ef
00
e6
00
00
00
01
01
00
00
00
02
00
fe
01
00
00
00
01
00
00
03
01
01
10
10
00
01
01
00
02
00
00
00
00
01
00
00
01
01
00
00
00
00
00
00
00
db
dd
fe
df
00
10
10
00
11
00
00
0b
dd
01
10
10
00
00
dc
d8
fe
dc
d9
01
10
10
00
11
00
00
00
00
00
00
00
00
00
00
04
d5
00
10
01
10
00
01
01
01
01
00
00
02
ce
00
00
00
00
f4
00
00
00
00
fa
