01
00
07
c4
80
87
46
07
87
00
f0
07
27
d6
f6
8a
07
a2
80
07
27
d7
8c
07
a5
75
80
01
24
20
26
22
04
09
24
09
94
20
f0
65
20
12
20
24
24
29
01
80
01
f7
26
24
22
20
2e
2c
2a
28
87
27
fe
07
a4
54
74
10
04
07
07
a8
27
99
84
f7
e7
20
09
89
0a
00
14
07
a0
07
16
07
87
07
a0
f0
a0
09
16
04
f0
19
09
0a
04
09
04
74
04
85
05
86
04
00
0a
89
1c
26
f7
87
27
07
fc
07
a8
07
80
04
04
0a
09
0a
20
f0
08
1a
07
20
f0
05
f0
05
f0
04
09
27
c2
05
f0
25
05
35
f0
20
f0
2b
f0
09
0b
00
84
f0
20
f0
05
f0
27
80
f0
07
27
45
75
15
f7
e7
20
80
07
a5
55
75
80
07
a5
15
55
80
07
a5
15
55
80
07
27
75
15
f7
e7
20
80
01
24
22
20
26
09
84
04
f0
1e
f0
08
07
07
a8
07
07
07
9e
f0
08
07
07
a8
05
f0
f0
1e
f0
f0
08
07
07
a8
07
07
07
92
f0
08
07
07
a8
20
24
24
29
01
80
06
c6
87
20
f0
26
86
87
80
f0
01
07
05
2e
24
f0
05
05
06
f0
05
f0
47
47
45
20
97
17
e7
e5
01
80
01
28
2e
2c
2a
26
09
17
f6
20
24
07
07
a8
24
29
29
01
80
07
07
80
d7
80
97
95
d5
d5
67
04
05
04
91
09
f0
f0
1e
f0
08
07
07
a8
07
07
07
e4
f0
08
07
07
a8
05
f0
f0
1e
f0
f0
08
07
07
a8
07
a7
87
00
a7
00
a7
00
a7
00
07
18
f0
0a
07
87
07
a0
24
20
24
29
29
05
01
f0
86
c6
87
20
f0
a6
06
07
80
f0
