// maybe we don't actually need it
module fpu(
    input opcode[6:0]


);


endmodule